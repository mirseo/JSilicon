// 헤드 연산 할당 장치

`define default_netname none

(* keep_hierarchy *)
module FSM(
    input wire clock,
    input wire reset,
    input wire tx
    );
endmodule