// 내부 레지스터 파일

`define default_netname none

(* keep_hierarchy *)
module REG (
    input wire clkm
    );
endmodule